//pack_top.v


module pack_top(



);



//---------------------------------------
//---------------------------------------



endmodule
