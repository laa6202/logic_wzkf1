//commu_m_push.v

module commu_m_push(

//clk rst
clk_sys,
rst_n
);

//clk rst
input clk_sys;
input rst_n;
//------------------------------------------
//------------------------------------------



endmodule
