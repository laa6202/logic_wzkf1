//syn_m_main.v

module syn_m_main(
fire_sync,
done_sync,
fire_info,
done_info,
//gps info
gps_pluse,
//clk rst
clk_sys,
pluse_us,
rst_n
);
output	fire_sync;
input		done_sync;
output	fire_info;
input		done_info;
//gps info
input		gps_pluse;
//clk rst
input clk_sys;
input pluse_us;
input rst_n;
//-------------------------------------------
//-------------------------------------------



endmodule
