//gps_source.v

module gps_source(
gps_pluse,
//clk rst
clk_sys,
rst_n
);
output gps_pluse;
//clk rst
input clk_sys;
input rst_n;
//-----------------------------------------
//-----------------------------------------


wire gps_pluse = 1'b0;


endmodule
