//commu_top.v

module commu_top(

//clk rst
clk_sys,
rst_n
);

//clk rst
input clk_sys;
input rst_n;
//--------------------------------------
//--------------------------------------



endmodule
