//commu_m_main.v

module commu_m_main(
fire_push,
done_push,
repk_frm,
buf_frm,
//configuration
arm_int_n,
stu_buf_rdy,
//clk rst
debug,
clk_sys,
rst_n
);
output	fire_push;
input		done_push;
input		repk_frm;
input 	buf_frm;
//configuration
output 	arm_int_n;
output [7:0] stu_buf_rdy;
//clk rst
output debug;
input clk_sys;
input rst_n;
//------------------------------------------
//------------------------------------------


reg repk_frm_reg;
reg buf_frm_reg;
always @(posedge clk_sys )	begin
	repk_frm_reg <= repk_frm;
	buf_frm_reg <= buf_frm;
end
wire repk_frm_falling = repk_frm_reg & (~repk_frm);
wire buf_frm_falling = buf_frm_reg & (~buf_frm);


reg arm_int;
always @(posedge clk_sys or negedge rst_n)	begin
	if(~rst_n)
		arm_int <= 1'b0;
	else if(buf_frm_falling)
		arm_int <= 1'b0;
	else if(repk_frm_falling)
		arm_int <= 1'b1;
	else ;
end

wire arm_int_n = ~arm_int;


wire [7:0] stu_buf_rdy;
assign stu_buf_rdy = arm_int_n ? 8'h0 : 8'hff;


//----------- for debug ------------
reg [9:0] cnt_repk_frm;
always @ (posedge clk_sys or negedge rst_n)	begin
	if(~rst_n)
		cnt_repk_frm <= 10'h0;
	else if(cnt_repk_frm  == 10'h3ff)
		;
	else if(buf_frm_falling)
		cnt_repk_frm <= cnt_repk_frm + 10'h1;
	else ;
end
wire debug = ^cnt_repk_frm;

endmodule
