//commu_m_top.v

module commu_m_top(
//arm spi
spi_csn,
spi_sck,
spi_miso,
spi_mosi,
//clk rst
clk_sys,
rst_n
);
input spi_csn;
input spi_sck;
output	spi_miso;
input		spi_mosi;

//clk rst
input clk_sys;
input rst_n;
//-----------------------------------------
//-----------------------------------------


endmodule
