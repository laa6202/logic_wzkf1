//commu_m_main.v

module commu_m_main(

//clk rst
clk_sys,
rst_n
);

//clk rst
input clk_sys;
input rst_n;
//------------------------------------------
//------------------------------------------



endmodule
