//syn_m_info.v

module syn_m_info(
tx_info,
fire_sync,
fire_info,
//clk rst
clk_sys,
rst_n
);

output	tx_info;
input		fire_sync;
input 	fire_info;
//clk rst
input clk_sys;
input rst_n;
//------------------------------------------
//------------------------------------------



endmodule

