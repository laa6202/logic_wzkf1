//fetch_top.v


module fetch_top(
rx_a,
rx_b,
//clk rst
fire_sync,
clk_sys,
rst_n
);

input rx_a;
input rx_b;
//clk rst
input fire_sync;
input clk_sys;
input rst_n;
//-----------------------------------------
//-----------------------------------------



endmodule

