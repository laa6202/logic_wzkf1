//commu_m_mux.v

module commu_m_mux(
req_rd,
req_q,
//configuratiuon
cfg_tp,
//clk rst
clk_sys,
rst_n
);
input					req_rd;
output [7:0]	req_q;
//configuratiuon
input [7:0]	cfg_tp;
//clk rst
input	clk_sys;
input rst_n;
//----------------------------------------
//----------------------------------------



endmodule
